BZh91AY&SY4z~� n߀py���߰����`<�l ��� @	����  �I4)驤       `��JT4&�22h ���� q�&LF& L�&@F ���D����     �F��i�M �4 �d��1D h�4Ѫ��ڈf��L�Hh6Bf���A
�T(|>!@��e~�����HMR�q�I$mDKm��!-��-�	e��B�^Y,��l���$'�B�;�E�D�H���O�y$�|���ň�0�A� �&�i���8to�����'䑤���S�J�H$ $	�8���A �A �H�*A"���$	����N	�"�8'��S�Z�	��(�$)kdV��	BT�pH'�H �B�i� �o�A �5)*�	�
�	�H ��d�D"��� �H���E%H4�H����x@g��Z��J������6���=�2"�=�쁇NvHt��X��Z�V�Bo.QA�64V]��K, �.v�ښ���mm�#/2Z6ʐn�̻�cԵ�ж̎�V�,c��a�m��n%`�P��h�æ¬��ib�.�R�-�6�b͞+��5�b��[��"�ke��^\Q�;J-u�Vػn[WF:4�:kˉ+�et�0�ƒ%�ն�[Ki��$���m��5ul���o����O��5���+(&+j�$��V�0q�TI!���%�n H����tJ��"�l�;���y~ztGF��j�q��&a�E �����	��Bb4{7p���eoRtR]�����u��m��6\t�O$���n��R�<s�n��ܝ{����Q�Ý�I��g8��{eq�e�:��"c�9)I$C%1B�8�;E{Y�0Xa3�A��n�C�uO�u��M$�ITtز(
�:�u�7vy���&J!�_d0.̂�~��v��X쪐
?B��k�XG8נ��Tss!�2����6��A���@ 4k��k�(�8Y*T�l����s�̔��_���������z�.���t�G����:������S�
. -{�1@;cB4
<��0S4Wu��Te?�x��j��JK��ȋ��?���{��=�eX��6�1�bfZhska��ݵ��Z�n l�%԰�����s�F1G�P�PF�J!�8�6U���@.�����o��g�YL���ExTM� .�>��q+~�a�%T�SiEA�u��/�<T
�� � :��X�!�:��h��,Zy�+O��妠�"�-v���$"�/|hp�zX��wLp��X�AF��M��L&A@H������{��.�(+(�x�x�#�
�׽�UURN�I'��l�����~�B���^uQ@��o�@>h�.���|(��=�pr�v�{���A)T�3U��^���s�i�+�=5�Y߄ j�Y�)á�G���L;�#;�� O:�l���4I�t� 9iT�E��]��i�i�'@�]���)IuB���Ba�Ǧ�ڬ�;"D��u�b%,��te��Z/���nJT�B�0��S�u_k����*�*͜5da��C�]W��o;�ʣ=A�6�
)�O���߹�$�]��Ӟ��x����-g	>+�~|8~���rTN��Q��
��%,H�7H�9;�C�jǆ�[=����s��O�e9�Y�f4+<>x�a�/��hp��N���f-�r���A=R�$$�ŌHڔ����
�θsCU-�Q�����*���5��� ��ڱl8��0�h����3��m���˿pw�ܿ@*�y$QF!���o�M=���8 ����g��t������yR�U*�*��QsUfy�4�:k�w|��xx�S�Y ���ʣ������
�p�r���ݤ�t��8�z��|m&^�=4kbs�˦)m�f���I�g��Ww��D�UPh`����x��}�x�E��}��:s�	s�L,#D��4S���I$*�9��B:�4�B:�� 0m�]�����1nM������e2���Uk�V�6L۹��3p±!����F�u���>�t@���(�C�=;Ӄ�����b�Y�mo���3Gw=H#�xzE�!A�C�k�������6��ʁ�Vt���(��=:��@�9��m���ԏ�r:���<�Q&�F��8�����Ă�"�:h��r��;�ןgX�1?J���a�<w���g���@g��=�9@x��x=���d yPW�F����v2$#'	#$�P
(� =+[�)�`ڬ��L���,ڮ�$\bZ+��T�KJp��
���
�	*�H��+j�&Pޖ��(-�� ��(���O�( �q�X /Z[ ri
����X����(�����kg��f�}F�����|A�s��'(��������Q��xx��R�'d��}n��=rBk(r��@�^��O����lK� ����9��3�ټB�|�F���s����qA� ~��J(_��!��u|d�&"PvG��~�y��ݶ�m��l��m��m��,�I!	$�I%|z3HE�fu��w�#M?��j��׎8����;��km��@��(i��)A��Q@�8E�n��X����;O��G�A�~���5  g��
 Kuƻ�C�r}Fߨ���׷�u6I��	�d_�ԟ8>�~.��"�S����������꛻@��;Jȭ����XP�ߡC�>��^F���n=������1�߬{DP�zd�����_�v+ ݬ8AQ������1MS�i�ò����y��ЧI`���:g��@ߦHo���87��P
V�>\��.$\K�Ԟ� `���a̽9\�*�h�  Z�p{��o�w�B(���W��i
�w_��yh��xG5�|�*��0��z�x���u����@j�� �M�;�<����@X���r4���>`�vb���J`��(�}W
���P�08q�;�tA՝����-���b­�㯯!	қSf0�U)�]���PV wl莇B9��r�Ӣw�(��8�}�&�O��8�'��l�î���H?��p��I��{�5f��]��B@����